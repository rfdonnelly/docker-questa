module hello_world;
initial $display("hello world");
endmodule
